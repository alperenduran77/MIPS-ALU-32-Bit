module xor_gate(
    input [31:0] a,
    input [31:0] b,
    output [31:0] y
);

    
    xor xor_gate_0(y[0], a[0], b[0]);
    xor xor_gate_1(y[1], a[1], b[1]);
	 xor xor_gate_2(y[2], a[2], b[2]);
	 xor xor_gate_3(y[3], a[3], b[3]);
	 xor xor_gate_4(y[4], a[4], b[4]);
	 xor xor_gate_5(y[5], a[5], b[5]);
	 xor xor_gate_6(y[6], a[6], b[6]);
	 xor xor_gate_7(y[7], a[7], b[7]);
	 xor xor_gate_8(y[8], a[8], b[8]);
	 xor xor_gate_9(y[9], a[9], b[9]);
	 xor xor_gate_10(y[10], a[10], b[10]);
    xor xor_gate_11(y[11], a[11], b[11]);
	 xor xor_gate_12(y[12], a[12], b[12]);
	 xor xor_gate_13(y[13], a[13], b[13]);
	 xor xor_gate_14(y[14], a[14], b[14]);
	 xor xor_gate_15(y[15], a[15], b[15]);
	 xor xor_gate_16(y[16], a[16], b[16]);
	 xor xor_gate_17(y[17], a[17], b[17]);
	 xor xor_gate_18(y[18], a[18], b[18]);
	 xor xor_gate_19(y[19], a[19], b[19]);
	 xor xor_gate_20(y[20], a[20], b[20]);
	 xor xor_gate_21(y[21], a[21], b[21]);
	 xor xor_gate_22(y[22], a[22], b[22]);
	 xor xor_gate_23(y[23], a[23], b[23]);
	 xor xor_gate_24(y[24], a[24], b[24]);
	 xor xor_gate_25(y[25], a[25], b[25]);
	 xor xor_gate_26(y[26], a[26], b[26]);
	 xor xor_gate_27(y[27], a[27], b[27]);
	 xor xor_gate_28(y[28], a[28], b[28]);
	 xor xor_gate_29(y[29], a[29], b[29]);
	 xor xor_gate_30(y[30], a[30], b[30]);
    xor xor_gate_31(y[31], a[31], b[31]);

endmodule
